LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL; 

PACKAGE mem_components IS

COMPONENT tri_buf
	GENERIC( N: INTEGER := 4);
	PORT ( 	X 	: IN STD_LOGIC_VECTOR (N-1 DOWNTO 0);
			E	: IN STD_LOGIC;
			F	: OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0 )); 
END COMPONENT; 

COMPONENT n_register
	GENERIC (N:INTEGER :=4);
	PORT (	R		:	IN	STD_LOGIC_VECTOR (N-1 DOWNTO 0);
			Rin,Clk	:	IN	STD_LOGIC; 
			Q		:	OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0)); 		
END COMPONENT; 

END mem_components; 

