LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL; 

ENTITY n_register IS
	GENERIC (N:INTEGER :=4);
	PORT (	R		:	IN	STD_LOGIC_VECTOR (N-1 DOWNTO 0);
			Rin,Clk	:	IN	STD_LOGIC; 
			Q		:	OUT STD_LOGIC_VECTOR (N-1 DOWNTO 0)); 
			
END n_register; 

ARCHITECTURE how_to_reg OF n_register IS 
BEGIN
	PROCESS (Clk)
	BEGIN
		IF RISING_EDGE (Clk) THEN
			IF Rin ='1' THEN
				Q<= R; 
			END IF; 
		END IF; 
	END PROCESS;
END how_to_reg; 